library verilog;
use verilog.vl_types.all;
entity aes_vlg_vec_tst is
end aes_vlg_vec_tst;
