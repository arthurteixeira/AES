library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity tb_top is
end entity;

architecture behavior of tb_top is


signal clock_sg     : std_logic := '0';
signal selInicio_sg : std_logic := '0';
signal selRound_sg  : std_logic := '0';
signal selKey_sg    : std_logic_vector(3 downto 0) := "0000";
signal enRegInicio_sg  : std_logic := '0';
signal enRegADR_sg     : std_logic := '0';
signal enRegSub_sg     : std_logic := '0';
signal enRegSR_sg      : std_logic := '0';
signal enRegMix_sg     : std_logic := '0';
signal enRegADR2_sg    : std_logic := '0';
signal plainText_sg : std_logic_vector(127 downto 0) := x"328831E0435A3137F6309807A88DA234";   -- (0 => '0', others=>'0');
signal keyIni_sg    : std_logic_vector(127 downto 0) :=   x"2B28AB097EAEF7CF15D2154F16A6883C"; -- (0 => '0', others=>'0');
signal outAes_sg    : std_logic_vector(127 downto 0);

component aes is
	port(
		clock                  : std_logic;
		selInicio 		 		  : std_logic;
		selRound               : std_logic;
		selKey                 : std_logic_vector(3 downto 0);
		enRegInicio            : std_logic;
		enRegADR               : std_logic;
		enRegSub               : std_logic;
		enRegSR                : std_logic;
		enRegMix               : std_logic;
		enRegADR2              : std_logic;
		plainText	           : in std_logic_vector(127 downto 0);
		keyIni     	           : in std_logic_vector(127 downto 0);
		outAes  : out std_logic_vector(127 downto 0)
	);
end component aes;

begin

inst_aes : aes
	port map(
		clock => clock_sg,
		selInicio => selInicio_sg,
		selRound => selRound_sg,
		selKey => selKey_sg,
		enRegInicio => enRegInicio_sg,
		enRegADR    => enRegADR_sg,
		enRegSub    => enRegSub_sg,        
		enRegSR     => enRegSR_sg,           
		enRegMix    => enRegMix_sg,           
		enRegADR2   => enRegADR2_sg,
		plainText => plainText_sg,
		keyIni => keyIni_sg,
		outAes => outAes_sg
	);
--lll
clock_sg <= not clock_sg after 20 ns;

process is
	begin			
		wait for 5 ns;
			enRegInicio_sg <= '1';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '0';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '1';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '0';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '1';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '0';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '1';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '0';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '1';           
			enRegADR2_sg   <= '0';
			selInicio_sg <= '1';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '1';
			selKey_sg         <= "0001";
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '1';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '0';
			selInicio_sg   <= '1';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '1';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '0';
			selInicio_sg   <= '0';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '1';           
			enRegADR2_sg   <= '0';
			selInicio_sg   <= '1';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '1';
			selInicio_sg   <= '0';
			selKey_sg         <= "0010";
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '1';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '0';
			selInicio_sg   <= '1';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '1';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '0';
			selInicio_sg   <= '0';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '1';           
			enRegADR2_sg   <= '0';
			selInicio_sg   <= '1';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '1';
			selInicio_sg   <= '0';
			selKey_sg         <= "0011";
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '1';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '0';
			selInicio_sg   <= '1';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '1';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '0';
			selInicio_sg   <= '0';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '1';           
			enRegADR2_sg   <= '0';
			selInicio_sg   <= '1';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '1';
			selInicio_sg   <= '0';
			selKey_sg         <= "0100";
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '1';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '0';
			selInicio_sg   <= '1';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '1';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '0';
			selInicio_sg   <= '0';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '1';           
			enRegADR2_sg   <= '0';
			selInicio_sg   <= '1';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '1';
			selInicio_sg   <= '0';
			selKey_sg         <= "0101";
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '1';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '0';
			selInicio_sg   <= '1';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '1';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '0';
			selInicio_sg   <= '0';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '1';           
			enRegADR2_sg   <= '0';
			selInicio_sg   <= '1';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '1';
			selInicio_sg   <= '0';
			selKey_sg         <= "0110";
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '1';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '0';
			selInicio_sg   <= '1';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '1';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '0';
			selInicio_sg   <= '0';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '1';           
			enRegADR2_sg   <= '0';
			selInicio_sg   <= '1';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '1';
			selInicio_sg   <= '0';
			selKey_sg         <= "0111";
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '1';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '0';
			selInicio_sg   <= '1';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '1';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '0';
			selInicio_sg   <= '0';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '1';           
			enRegADR2_sg   <= '0';
			selInicio_sg   <= '1';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '1';
			selInicio_sg   <= '0';
			selKey_sg         <= "1000";
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '1';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '0';
			selInicio_sg   <= '1';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '1';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '0';
			selInicio_sg   <= '0';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '1';           
			enRegADR2_sg   <= '0';
			selInicio_sg   <= '1';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '1';
			selInicio_sg   <= '0';
			selKey_sg         <= "1001";
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '1';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '0';
			selInicio_sg   <= '1';
			selRound_sg    <= '1';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '1';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '0';
			selInicio_sg   <= '0';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '1';           
			enRegADR2_sg   <= '0';
			selInicio_sg   <= '1';
		wait for 40 ns;
			enRegInicio_sg <= '0';
			enRegADR_sg    <= '0';
			enRegSub_sg    <= '0';           
			enRegSR_sg     <= '0';           
			enRegMix_sg    <= '0';           
			enRegADR2_sg   <= '1';
			selInicio_sg   <= '0';
			selKey_sg         <= "1010";
		wait;	
end process;
	
end behavior;

